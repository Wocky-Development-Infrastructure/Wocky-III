module wockyfx

import core.wocky

pub struct WockyFX {

}