/*
	List of online users
*/
module commands