module scanner

