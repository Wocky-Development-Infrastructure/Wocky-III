module wocky