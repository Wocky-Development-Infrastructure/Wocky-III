/*	
	List of online bots
*/
module commands