module commands