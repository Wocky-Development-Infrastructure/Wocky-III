module thread_system

pub struct Threads {
	pub mut:
		thread_id		int
}