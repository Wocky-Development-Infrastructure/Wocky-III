module tools

import os
import net.http

pub fn geoip() {

}

pub fn dblookup() {

}

pub fn cfresolver() {
	
}
