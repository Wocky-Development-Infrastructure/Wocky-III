module term_control


// Return a string with the color in ANSI Escape sequence code
pub fn rgb_ansi(rgb []string) string {
	return ""
}