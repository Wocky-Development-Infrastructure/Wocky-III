module crud

import os
import mysql

pub fn create_api(api string, mut sql mysql.Connection)  {

}

pub fn read_api(api string, mut sql mysql.Connection)  {

}

pub fn update_api(api string, mut sql mysql.Connection)  {

}

pub fn delete_api(api string, mut sql mysql.Connection)  {

}