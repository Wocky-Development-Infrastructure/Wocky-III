/*
	User must confirm the current password
*/
module commands