module crud

import os
import mysql
