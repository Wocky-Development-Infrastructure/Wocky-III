module term_control

pub fn gradiant(startrgb, endrgb, text) {

}
