module logger

pub fn send_error() {

}

pub fn send_cmd_log() {

}

pub fn send_login_log() {

}

pub fn send_attack_log() {

}

pub fn send_admin_log() {

}